module clap

pub struct Command {
pub:
	name string [required]
	description string
}