module clap

pub struct Flag {
pub mut:
	value int
}