// module main

// import clap

// fn main() {
// 	flag := clap.Flag{name: 'test'}
// 	println(flag.name)
// }
